
module SevenSegment(


	output		     [7:0]		hex,
	input 		     [3:0]		bin,
	input 		     				point
);
reg [6:0] led;
assign hex[6:0]=~led[6:0];
assign hex[7] = ~point;
//sets up a reg for the seven segment display
//inverts all data so that it turns on the proper parts of the display

always @ (bin[3:0]) begin//case statement that turns on the proper parts of the seven segment led for the corresponding number
case(bin[3:0])
4'b0000:begin
led[0]=1;
led[1]=1;
led[2]=1;
led[3]=1;
led[4]=1;
led[5]=1;
led[6]=0;
end
4'b0001:begin
led[0]=0;
led[1]=1;
led[2]=1;
led[3]=0;
led[4]=0;
led[5]=0;
led[6]=0;
end
4'b0010:begin
led[0]=1;
led[1]=1;
led[2]=0;
led[3]=1;
led[4]=1;
led[5]=0;
led[6]=1;
end
4'b0011:begin
led[0]=1;
led[1]=1;
led[2]=1;
led[3]=1;
led[4]=0;
led[5]=0;
led[6]=1;
end
4'b0100:begin
led[0]=0;
led[1]=1;
led[2]=1;
led[3]=0;
led[4]=0;
led[5]=1;
led[6]=1;
end
4'b0101:begin
led[0]=1;
led[1]=0;
led[2]=1;
led[3]=1;
led[4]=0;
led[5]=1;
led[6]=1;
end
4'b0110:begin
led[0]=1;
led[1]=0;
led[2]=1;
led[3]=1;
led[4]=1;
led[5]=1;
led[6]=1;
end
4'b0111:begin
led[0]=1;
led[1]=1;
led[2]=1;
led[3]=0;
led[4]=0;
led[5]=0;
led[6]=0;
end
4'b1000:begin
led[0]=1;
led[1]=1;
led[2]=1;
led[3]=1;
led[4]=1;
led[5]=1;
led[6]=1;
end
4'b1001:begin
led[0]=1;
led[1]=1;
led[2]=1;
led[3]=0;
led[4]=0;
led[5]=1;
led[6]=1;
end
4'b1010:begin
led[0]=1;
led[1]=1;
led[2]=1;
led[3]=0;
led[4]=1;
led[5]=1;
led[6]=1;
end
4'b1011:begin
led[0]=0;
led[1]=0;
led[2]=1;
led[3]=1;
led[4]=1;
led[5]=1;
led[6]=1;
end
4'b1100:begin
led[0]=1;
led[1]=0;
led[2]=0;
led[3]=1;
led[4]=1;
led[5]=1;
led[6]=0;
end
4'b1101:begin
led[0]=0;
led[1]=1;
led[2]=1;
led[3]=1;
led[4]=1;
led[5]=0;
led[6]=1;
end
4'b1110:begin
led[0]=1;
led[1]=0;
led[2]=0;
led[3]=1;
led[4]=1;
led[5]=1;
led[6]=1;
end
4'b1111:begin
led[0]=1;
led[1]=0;
led[2]=0;
led[3]=0;
led[4]=1;
led[5]=1;
led[6]=1;
end
default:begin
led[0]=0;
led[1]=0;
led[2]=0;
led[3]=0;
led[4]=0;
led[5]=0;
led[6]=0;
end
endcase
end
endmodule
